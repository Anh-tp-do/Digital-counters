// Ring counter 

module ring_counter(d, clk, out);
  input d, clk;
  output out;
  
  always @(posedge clk)
    begin
      if (!rst)
        
    end 
endmodule 
